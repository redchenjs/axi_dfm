/*
 * config.sv
 *
 *  Created on: 2021-05-21 19:25
 *      Author: Jack Chen <redchenjs@live.com>
 */

parameter [32:0] DEFAULT_GATE_TIME = 32'd24_999;
