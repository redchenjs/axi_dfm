/*
 * config.sv
 *
 *  Created on: 2021-05-21 19:25
 *      Author: Jack Chen <redchenjs@live.com>
 */

parameter [3:0] RTL_REVISION_MAJOR = 4'h1;
parameter [3:0] RTL_REVISION_MINOR = 4'h0;

parameter [32:0] DEFAULT_GATE_TIME = 32'd199_999;
