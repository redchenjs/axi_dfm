/*
 * test_ram_rw.sv
 *
 *  Created on: 2020-07-19 18:00
 *      Author: Jack Chen <redchenjs@live.com>
 */

`timescale 1ns / 1ps

module test_measure;

logic clk_i;
logic rst_n_i;

logic sig_clk_i;

logic [5:0] ref_clk_i;
logic [5:0] ref_rst_n_i;

logic        reg_wr_en_o;
logic [63:0] reg_wr_data_o;

measure measure(
    .clk_i(clk_i),
    .rst_n_i(rst_n_i),

    .sig_clk_i(sig_clk_i),

    .ref_clk_i(ref_clk_i),
    .ref_rst_n_i(ref_rst_n_i),

    .reg_wr_en_o(reg_wr_en_o),
    .reg_wr_data_o(reg_wr_data_o)
);

initial begin
    clk_i   <= 1'b1;
    rst_n_i <= 1'b0;

    sig_clk_i <= 1'b1;

    ref_clk_i   <= 6'h00;
    ref_rst_n_i <= 6'h00;

    #2 rst_n_i <= 1'b1;
    #2 ref_rst_n_i <= 6'h3f;
end

always begin
    #2.4 clk_i <= ~clk_i;
end

always begin
    #250 sig_clk_i <= ~sig_clk_i;
end

always begin
    while (1) begin
        #2.4 ref_clk_i[0] <= ~ref_clk_i[0];
    end
end

always begin
    #0.8
    while (1) begin
        #2.4 ref_clk_i[1] <= ~ref_clk_i[1];
    end
end

always begin
    #1.6
    while (1) begin
        #2.4 ref_clk_i[2] <= ~ref_clk_i[2];
    end
end

always begin
    #2.4
    while (1) begin
        #2.4 ref_clk_i[3] <= ~ref_clk_i[3];
    end
end

always begin
    #3.2
    while (1) begin
        #2.4 ref_clk_i[4] <= ~ref_clk_i[4];
    end
end

always begin
    #4.0
    while (1) begin
        #2.4 ref_clk_i[5] <= ~ref_clk_i[5];
    end
end

always begin
    #1000000 rst_n_i <= 1'b0;

    #25 $stop;
end

endmodule
