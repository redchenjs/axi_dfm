/*
 * config.sv
 *
 *  Created on: 2021-05-21 19:25
 *      Author: Jack Chen <redchenjs@live.com>
 */

`ifndef _CONFIG_SV_
`define _CONFIG_SV_

localparam [31:0] DEFAULT_GATE_TIME_SHIFT = 32'd49_999;
localparam [31:0] DEFAULT_GATE_TIME_TOTAL = 32'd249_999;

`endif
